class uart_monitor extends uvm_component;

endclass