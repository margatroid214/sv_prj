class apb_base_seq extends uvm_sequence #(apb_seq_item);
  function new
endclass