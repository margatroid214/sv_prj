`include "uvm_pkg.sv"

package apbuart_env_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import uart_cfg_pkg::*;
import apb_agent_pkg::*;
import uart_agent_pkg::*;

`include "../config/apbuart_macros.sv"
//`include "../agents/apb_agent/apb_if.sv"
//`include "../agents/uart_agent/uart_if.sv"

`include "vsequencer.sv"
`include "apb_seq_lib.sv"
`include "uart_seq_lib.sv"
`include "apbuart_vseq_lib.sv"
`include "apbuart_model.sv"
`include "apbuart_scoreboard.sv"
`include "apbuart_env.sv"
`include "apbuart_test_lib.sv"

endpackage