class apbuart_env extends uvm_env;

endclass