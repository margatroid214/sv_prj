
package apb_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "apb_seq_item.sv"

endpackage