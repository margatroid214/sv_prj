package uart_agent_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "uart_transaction.sv"

endpackage