class apb_cov extends uvm_subscriber #(apb_seq_item);

endclass